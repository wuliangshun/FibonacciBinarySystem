module RAM_fibonacci(rst,cnt_a,mema);
input rst;
input [9:0] cnt_a;
output reg [15:0] mema;
 reg  [63:0] mem[127:0];
  always@(negedge rst) begin 
        mem[0]=0;
mem[1]=1;
mem[2]=1;
mem[3]=2;
mem[4]=3;
mem[5]=5;
mem[6]=8;
mem[7]=13;
mem[8]=21;
mem[9]=34;
mem[10]=55;
mem[11]=89;
mem[12]=144;
mem[13]=233;
mem[14]=377;
mem[15]=610;
mem[16]=987;
mem[17]=1597;
mem[18]=2584;
mem[19]=4181;
mem[20]=6765;
mem[21]=10946;
mem[22]=17711;
mem[23]=28657;
mem[24]=46368;
mem[25]=75025;
mem[26]=121393;
mem[27]=196418;
mem[28]=317811;
mem[29]=514229;
mem[30]=832040;
mem[31]=1346269;
mem[32]=2178309;
mem[33]=3524578;
mem[34]=5702887;
mem[35]=9227465;
mem[36]=14930352;
mem[37]=24157817;
mem[38]=39088169;
mem[39]=63245986;
mem[40]=102334155;
mem[41]=165580141;
mem[42]=267914296;
mem[43]=433494437;
mem[44]=701408733;
mem[45]=1134903170;
mem[46]=1836311903;
mem[47]=2971215073;
mem[48]=4807526976;
mem[49]=7778742049;
mem[50]=12586269025;
mem[51]=20365011074;
mem[52]=32951280099;
mem[53]=53316291173;
mem[54]=86267571272;
mem[55]=139583862445;
mem[56]=225851433717;
mem[57]=365435296162;
mem[58]=591286729879;
mem[59]=956722026041;
mem[60]=1548008755920;
mem[61]=2504730781961;
mem[62]=4052739537881;
mem[63]=6557470319842;
mem[64]=10610209857723;
mem[65]=17167680177565;
mem[66]=27777890035288;
mem[67]=44945570212853;
mem[68]=72723460248141;
mem[69]=117669030460994;
mem[70]=190392490709135;
mem[71]=308061521170129;
mem[72]=498454011879264;
mem[73]=806515533049393;
mem[74]=1304969544928657;
mem[75]=2111485077978050;
mem[76]=3416454622906707;
mem[77]=5527939700884757;
mem[78]=8944394323791464;
mem[79]=14472334024676221;
mem[80]=23416728348467685;
mem[81]=37889062373143906;
mem[82]=61305790721611591;
mem[83]=99194853094755497;
mem[84]=160500643816367088;
mem[85]=259695496911122585;
mem[86]=420196140727489673;
mem[87]=679891637638612258;
mem[88]=1100087778366101931;
mem[89]=1779979416004714189;
mem[90]=2880067194370816120;
mem[91]=4660046610375530309;
mem[92]=7540113804746346429;
mem[93]=12200160415121876738;
mem[94]=19740274219868223167;
mem[95]=31940434634990099905;
mem[96]=51680708854858323072;
mem[97]=83621143489848422977;
mem[98]=135301852344706746049;
mem[99]=218922995834555169026;
mem[100]=354224848179261915075;
mem[101]=573147844013817084101;
mem[102]=927372692193078999176;
mem[103]=1500520536206896083277;
mem[104]=2427893228399975082453;
mem[105]=3928413764606871165730;
mem[106]=6356306993006846248183;
mem[107]=10284720757613717413913;
mem[108]=16641027750620563662096;
mem[109]=26925748508234281076009;
mem[110]=43566776258854844738105;
mem[111]=70492524767089125814114;
mem[112]=114059301025943970552219;
mem[113]=184551825793033096366333;
mem[114]=298611126818977066918552;
mem[115]=483162952612010163284885;
mem[116]=781774079430987230203437;
mem[117]=1264937032042997393488322;
mem[118]=2046711111473984623691759;
mem[119]=3311648143516982017180081;
mem[120]=5358359254990966640871840;
mem[121]=8670007398507948658051921;
mem[122]=14028366653498915298923761;
mem[123]=22698374052006863956975682;
mem[124]=36726740705505779255899443;
mem[125]=59425114757512643212875125;
mem[126]=96151855463018422468774568;
mem[127]=155576970220531065681649693;
    end 
	 always@(cnt_a)begin
	     mema=mem[cnt_a];
	 end 
endmodule  
